`ifndef CFS_ALGN_PKG_SV
`define CFS_ALGN_PKG_SV

package cfs_algn_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "cfs_algn_env.sv"

endpackage

`endif
