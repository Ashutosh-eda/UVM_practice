`ifndef CFS_APB_TYPES_SV
  `define CFS_APB_TYPES_SV

    //Virtual interface type
    typedef virtual cfs_apb_if cfs_apb_vif;

`endif
